localparam[BYTE_WIDTH-1:0]
  F9PCAP_SEQNO_LENGTH     = 4,
  RECOVER_REQ_COUNT_L     = 2, // RecoverCount
  RECOVER_REQ_ADDR_FROM_L = 4, // AddrFrom
  RECOVER_REQ_ADDR_FROM_W = RECOVER_REQ_ADDR_FROM_L * BYTE_WIDTH,
  RECOVER_REQ_CHECK_L     = 8, // CheckData = [TTL]
  RECOVER_REQ_LENGTH = F9PCAP_SEQNO_LENGTH + RECOVER_REQ_COUNT_L + RECOVER_REQ_ADDR_FROM_L + RECOVER_REQ_CHECK_L,

  RECOVER_REQ_WIDTH  = RECOVER_REQ_LENGTH  * BYTE_WIDTH,
  F9PCAP_SEQNO_WIDTH = F9PCAP_SEQNO_LENGTH * BYTE_WIDTH,

  F9PCAP_EXT_HDR_LENGTH = F9PCAP_SEQNO_LENGTH + RECOVER_REQ_ADDR_FROM_L,
  F9PCAP_EXT_HDR_WIDTH  = F9PCAP_EXT_HDR_LENGTH * BYTE_WIDTH,

  // last_seqno             [F9PCAP_SEQNO_LENGTH    ]
  // last_addr              [RECOVER_REQ_ADDR_FROM_L]
  // last_recover_req_seqno [F9PCAP_SEQNO_LENGTH    ]
  // last_recover_req_addr  [RECOVER_REQ_ADDR_FROM_L]
  // last_recover_result    [ 1]
  DEV_ST_RECOVER_INFO_L = F9PCAP_SEQNO_LENGTH*2 + RECOVER_REQ_ADDR_FROM_L*2 + 1,
  DEV_ST_RECOVER_INFO_W = DEV_ST_RECOVER_INFO_L * BYTE_WIDTH,
